module tb_top_axi_serdes;

// Make sure to call finish so test exits
always begin
    $finish();
end

endmodule