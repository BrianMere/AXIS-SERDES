module top_axi_serdes(
    input clk
);

    // Start coding here... 

endmodule 